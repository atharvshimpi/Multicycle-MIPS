/*##########################################################################################
Note: Please don’t upload the assignments, template file/solution and lab. manual on GitHub or others public repository. 
Kindly remove them, if you have uploaded the previous assignments. 
It violates the BITS’s Intellectual Property Rights (IPR).
*******************************************************************************************/


module forwardingUnit(input [4:0] rs_id, input [4:0] rt_id, input [4:0] rs_ex, input [4:0] rt_ex, input [4:0] rd_mem, 
                        input [4:0] rd_wb, input regwrite_mem, input regwrite_wb, 
                        output reg [1:0] forward_a, output reg [1:0] forward_b, output reg forward_c, output reg forward_ad, output reg forward_bd);
    
    //WRITE YOUR CODE HERE
    

endmodule

